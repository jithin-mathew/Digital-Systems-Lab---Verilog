module full_adder(a,b,cin,sum,cout);
input a;
input b;
input cin;
output sum;
output cout;

assign sum = a^b^cin;
assign cout = (a & b) | (cin & (a^b)); 

endmodule

module bitadder(A,B,Cin,Sum,Cout);

input [3:0]A;
input [3:0]B;
input Cin;

output [3:0]Sum;
output Cout;

wire c1,c2,c3;

full_adder f1(.a(A[0]),.b(B[0]),.cin(Cin),.sum(Sum[0]),.cout(c1));
full_adder f2(.a(A[1]),.b(B[1]),.cin(c1),.sum(Sum[1]),.cout(c2));
full_adder f3(.a(A[2]),.b(B[2]),.cin(c2),.sum(Sum[2]),.cout(c3));
full_adder f4(.a(A[3]),.b(B[3]),.cin(c3),.sum(Sum[3]),.cout(Cout));

endmodule

module testbench();
reg [3:0]A;
reg [3:0]B;
reg Cin;
wire [3:0]Sum;
wire Cout;

bitadder tb(A,B,Cin,Sum,Cout);

initial
begin

$monitor("A = %b : B = %b : Cin = %b : Sum = %b : Cout = %b ",A,B,Cin,Sum,Cout);
$dumpfile("4bitadder.vcd");
$dumpvars;

A = 4'b0000 ; B = 4'b0000 ; Cin = 1'b0 ;
#5; 
A = 4'b0000 ; B = 4'b0001 ; Cin = 1'b0 ;
#5; 
A = 4'b0000 ; B = 4'b0010 ; Cin = 1'b0 ;
#5; 
A = 4'b0000 ; B = 4'b0011 ; Cin = 1'b0 ;
#5; 
A = 4'b0000 ; B = 4'b0100 ; Cin = 1'b0 ;
#5; 
A = 4'b0000 ; B = 4'b0101 ; Cin = 1'b0 ;
#5; 
A = 4'b0000 ; B = 4'b0110 ; Cin = 1'b0 ;
#5; 
A = 4'b0000 ; B = 4'b0111 ; Cin = 1'b0 ;
#5; 
A = 4'b0000 ; B = 4'b1000 ; Cin = 1'b0 ;
#5; 
A = 4'b0000 ; B = 4'b1001 ; Cin = 1'b0 ;
#5; 
A = 4'b0000 ; B = 4'b1010 ; Cin = 1'b0 ;
#5; 
A = 4'b0000 ; B = 4'b1011 ; Cin = 1'b0 ;
#5; 
A = 4'b0000 ; B = 4'b1100 ; Cin = 1'b0 ;
#5; 
A = 4'b0000 ; B = 4'b1101 ; Cin = 1'b0 ;
#5; 
A = 4'b0000 ; B = 4'b1110 ; Cin = 1'b0 ;
#5; 
A = 4'b0000 ; B = 4'b1111 ; Cin = 1'b0 ;
#5; 
A = 4'b0001 ; B = 4'b0000 ; Cin = 1'b0 ;
#5; 
A = 4'b0001 ; B = 4'b0001 ; Cin = 1'b0 ;
#5; 
A = 4'b0001 ; B = 4'b0010 ; Cin = 1'b0 ;
#5; 
A = 4'b0001 ; B = 4'b0011 ; Cin = 1'b0 ;
#5; 
A = 4'b0001 ; B = 4'b0100 ; Cin = 1'b0 ;
#5; 
A = 4'b0001 ; B = 4'b0101 ; Cin = 1'b0 ;
#5; 
A = 4'b0001 ; B = 4'b0110 ; Cin = 1'b0 ;
#5; 
A = 4'b0001 ; B = 4'b0111 ; Cin = 1'b0 ;
#5; 
A = 4'b0001 ; B = 4'b1000 ; Cin = 1'b0 ;
#5; 
A = 4'b0001 ; B = 4'b1001 ; Cin = 1'b0 ;
#5; 
A = 4'b0001 ; B = 4'b1010 ; Cin = 1'b0 ;
#5; 
A = 4'b0001 ; B = 4'b1011 ; Cin = 1'b0 ;
#5; 
A = 4'b0001 ; B = 4'b1100 ; Cin = 1'b0 ;
#5; 
A = 4'b0001 ; B = 4'b1101 ; Cin = 1'b0 ;
#5; 
A = 4'b0001 ; B = 4'b1110 ; Cin = 1'b0 ;
#5; 
A = 4'b0001 ; B = 4'b1111 ; Cin = 1'b0 ;
#5; 
A = 4'b0010 ; B = 4'b0000 ; Cin = 1'b0 ;
#5; 
A = 4'b0010 ; B = 4'b0001 ; Cin = 1'b0 ;
#5; 
A = 4'b0010 ; B = 4'b0010 ; Cin = 1'b0 ;
#5; 
A = 4'b0010 ; B = 4'b0011 ; Cin = 1'b0 ;
#5; 
A = 4'b0010 ; B = 4'b0100 ; Cin = 1'b0 ;
#5; 
A = 4'b0010 ; B = 4'b0101 ; Cin = 1'b0 ;
#5; 
A = 4'b0010 ; B = 4'b0110 ; Cin = 1'b0 ;
#5; 
A = 4'b0010 ; B = 4'b0111 ; Cin = 1'b0 ;
#5; 
A = 4'b0010 ; B = 4'b1000 ; Cin = 1'b0 ;
#5; 
A = 4'b0010 ; B = 4'b1001 ; Cin = 1'b0 ;
#5; 
A = 4'b0010 ; B = 4'b1010 ; Cin = 1'b0 ;
#5; 
A = 4'b0010 ; B = 4'b1011 ; Cin = 1'b0 ;
#5; 
A = 4'b0010 ; B = 4'b1100 ; Cin = 1'b0 ;
#5; 
A = 4'b0010 ; B = 4'b1101 ; Cin = 1'b0 ;
#5; 
A = 4'b0010 ; B = 4'b1110 ; Cin = 1'b0 ;
#5; 
A = 4'b0010 ; B = 4'b1111 ; Cin = 1'b0 ;
#5; 
A = 4'b0011 ; B = 4'b0000 ; Cin = 1'b0 ;
#5; 
A = 4'b0011 ; B = 4'b0001 ; Cin = 1'b0 ;
#5; 
A = 4'b0011 ; B = 4'b0010 ; Cin = 1'b0 ;
#5; 
A = 4'b0011 ; B = 4'b0011 ; Cin = 1'b0 ;
#5; 
A = 4'b0011 ; B = 4'b0100 ; Cin = 1'b0 ;
#5; 
A = 4'b0011 ; B = 4'b0101 ; Cin = 1'b0 ;
#5; 
A = 4'b0011 ; B = 4'b0110 ; Cin = 1'b0 ;
#5; 
A = 4'b0011 ; B = 4'b0111 ; Cin = 1'b0 ;
#5; 
A = 4'b0011 ; B = 4'b1000 ; Cin = 1'b0 ;
#5; 
A = 4'b0011 ; B = 4'b1001 ; Cin = 1'b0 ;
#5; 
A = 4'b0011 ; B = 4'b1010 ; Cin = 1'b0 ;
#5; 
A = 4'b0011 ; B = 4'b1011 ; Cin = 1'b0 ;
#5; 
A = 4'b0011 ; B = 4'b1100 ; Cin = 1'b0 ;
#5; 
A = 4'b0011 ; B = 4'b1101 ; Cin = 1'b0 ;
#5; 
A = 4'b0011 ; B = 4'b1110 ; Cin = 1'b0 ;
#5; 
A = 4'b0011 ; B = 4'b1111 ; Cin = 1'b0 ;
#5; 
A = 4'b0100 ; B = 4'b0000 ; Cin = 1'b0 ;
#5; 
A = 4'b0100 ; B = 4'b0001 ; Cin = 1'b0 ;
#5; 
A = 4'b0100 ; B = 4'b0010 ; Cin = 1'b0 ;
#5; 
A = 4'b0100 ; B = 4'b0011 ; Cin = 1'b0 ;
#5; 
A = 4'b0100 ; B = 4'b0100 ; Cin = 1'b0 ;
#5; 
A = 4'b0100 ; B = 4'b0101 ; Cin = 1'b0 ;
#5; 
A = 4'b0100 ; B = 4'b0110 ; Cin = 1'b0 ;
#5; 
A = 4'b0100 ; B = 4'b0111 ; Cin = 1'b0 ;
#5; 
A = 4'b0100 ; B = 4'b1000 ; Cin = 1'b0 ;
#5; 
A = 4'b0100 ; B = 4'b1001 ; Cin = 1'b0 ;
#5; 
A = 4'b0100 ; B = 4'b1010 ; Cin = 1'b0 ;
#5; 
A = 4'b0100 ; B = 4'b1011 ; Cin = 1'b0 ;
#5; 
A = 4'b0100 ; B = 4'b1100 ; Cin = 1'b0 ;
#5; 
A = 4'b0100 ; B = 4'b1101 ; Cin = 1'b0 ;
#5; 
A = 4'b0100 ; B = 4'b1110 ; Cin = 1'b0 ;
#5; 
A = 4'b0100 ; B = 4'b1111 ; Cin = 1'b0 ;
#5; 
A = 4'b0101 ; B = 4'b0000 ; Cin = 1'b0 ;
#5; 
A = 4'b0101 ; B = 4'b0001 ; Cin = 1'b0 ;
#5; 
A = 4'b0101 ; B = 4'b0010 ; Cin = 1'b0 ;
#5; 
A = 4'b0101 ; B = 4'b0011 ; Cin = 1'b0 ;
#5; 
A = 4'b0101 ; B = 4'b0100 ; Cin = 1'b0 ;
#5; 
A = 4'b0101 ; B = 4'b0101 ; Cin = 1'b0 ;
#5; 
A = 4'b0101 ; B = 4'b0110 ; Cin = 1'b0 ;
#5; 
A = 4'b0101 ; B = 4'b0111 ; Cin = 1'b0 ;
#5; 
A = 4'b0101 ; B = 4'b1000 ; Cin = 1'b0 ;
#5; 
A = 4'b0101 ; B = 4'b1001 ; Cin = 1'b0 ;
#5; 
A = 4'b0101 ; B = 4'b1010 ; Cin = 1'b0 ;
#5; 
A = 4'b0101 ; B = 4'b1011 ; Cin = 1'b0 ;
#5; 
A = 4'b0101 ; B = 4'b1100 ; Cin = 1'b0 ;
#5; 
A = 4'b0101 ; B = 4'b1101 ; Cin = 1'b0 ;
#5; 
A = 4'b0101 ; B = 4'b1110 ; Cin = 1'b0 ;
#5; 
A = 4'b0101 ; B = 4'b1111 ; Cin = 1'b0 ;
#5; 
A = 4'b0110 ; B = 4'b0000 ; Cin = 1'b0 ;
#5; 
A = 4'b0110 ; B = 4'b0001 ; Cin = 1'b0 ;
#5; 
A = 4'b0110 ; B = 4'b0010 ; Cin = 1'b0 ;
#5; 
A = 4'b0110 ; B = 4'b0011 ; Cin = 1'b0 ;
#5; 
A = 4'b0110 ; B = 4'b0100 ; Cin = 1'b0 ;
#5; 
A = 4'b0110 ; B = 4'b0101 ; Cin = 1'b0 ;
#5; 
A = 4'b0110 ; B = 4'b0110 ; Cin = 1'b0 ;
#5; 
A = 4'b0110 ; B = 4'b0111 ; Cin = 1'b0 ;
#5; 
A = 4'b0110 ; B = 4'b1000 ; Cin = 1'b0 ;
#5; 
A = 4'b0110 ; B = 4'b1001 ; Cin = 1'b0 ;
#5; 
A = 4'b0110 ; B = 4'b1010 ; Cin = 1'b0 ;
#5; 
A = 4'b0110 ; B = 4'b1011 ; Cin = 1'b0 ;
#5; 
A = 4'b0110 ; B = 4'b1100 ; Cin = 1'b0 ;
#5; 
A = 4'b0110 ; B = 4'b1101 ; Cin = 1'b0 ;
#5; 
A = 4'b0110 ; B = 4'b1110 ; Cin = 1'b0 ;
#5; 
A = 4'b0110 ; B = 4'b1111 ; Cin = 1'b0 ;
#5; 
A = 4'b0111 ; B = 4'b0000 ; Cin = 1'b0 ;
#5; 
A = 4'b0111 ; B = 4'b0001 ; Cin = 1'b0 ;
#5; 
A = 4'b0111 ; B = 4'b0010 ; Cin = 1'b0 ;
#5; 
A = 4'b0111 ; B = 4'b0011 ; Cin = 1'b0 ;
#5; 
A = 4'b0111 ; B = 4'b0100 ; Cin = 1'b0 ;
#5; 
A = 4'b0111 ; B = 4'b0101 ; Cin = 1'b0 ;
#5; 
A = 4'b0111 ; B = 4'b0110 ; Cin = 1'b0 ;
#5; 
A = 4'b0111 ; B = 4'b0111 ; Cin = 1'b0 ;
#5; 
A = 4'b0111 ; B = 4'b1000 ; Cin = 1'b0 ;
#5; 
A = 4'b0111 ; B = 4'b1001 ; Cin = 1'b0 ;
#5; 
A = 4'b0111 ; B = 4'b1010 ; Cin = 1'b0 ;
#5; 
A = 4'b0111 ; B = 4'b1011 ; Cin = 1'b0 ;
#5; 
A = 4'b0111 ; B = 4'b1100 ; Cin = 1'b0 ;
#5; 
A = 4'b0111 ; B = 4'b1101 ; Cin = 1'b0 ;
#5; 
A = 4'b0111 ; B = 4'b1110 ; Cin = 1'b0 ;
#5; 
A = 4'b0111 ; B = 4'b1111 ; Cin = 1'b0 ;
#5; 
A = 4'b1000 ; B = 4'b0000 ; Cin = 1'b0 ;
#5; 
A = 4'b1000 ; B = 4'b0001 ; Cin = 1'b0 ;
#5; 
A = 4'b1000 ; B = 4'b0010 ; Cin = 1'b0 ;
#5; 
A = 4'b1000 ; B = 4'b0011 ; Cin = 1'b0 ;
#5; 
A = 4'b1000 ; B = 4'b0100 ; Cin = 1'b0 ;
#5; 
A = 4'b1000 ; B = 4'b0101 ; Cin = 1'b0 ;
#5; 
A = 4'b1000 ; B = 4'b0110 ; Cin = 1'b0 ;
#5; 
A = 4'b1000 ; B = 4'b0111 ; Cin = 1'b0 ;
#5; 
A = 4'b1000 ; B = 4'b1000 ; Cin = 1'b0 ;
#5; 
A = 4'b1000 ; B = 4'b1001 ; Cin = 1'b0 ;
#5; 
A = 4'b1000 ; B = 4'b1010 ; Cin = 1'b0 ;
#5; 
A = 4'b1000 ; B = 4'b1011 ; Cin = 1'b0 ;
#5; 
A = 4'b1000 ; B = 4'b1100 ; Cin = 1'b0 ;
#5; 
A = 4'b1000 ; B = 4'b1101 ; Cin = 1'b0 ;
#5; 
A = 4'b1000 ; B = 4'b1110 ; Cin = 1'b0 ;
#5; 
A = 4'b1000 ; B = 4'b1111 ; Cin = 1'b0 ;
#5; 
A = 4'b1001 ; B = 4'b0000 ; Cin = 1'b0 ;
#5; 
A = 4'b1001 ; B = 4'b0001 ; Cin = 1'b0 ;
#5; 
A = 4'b1001 ; B = 4'b0010 ; Cin = 1'b0 ;
#5; 
A = 4'b1001 ; B = 4'b0011 ; Cin = 1'b0 ;
#5; 
A = 4'b1001 ; B = 4'b0100 ; Cin = 1'b0 ;
#5; 
A = 4'b1001 ; B = 4'b0101 ; Cin = 1'b0 ;
#5; 
A = 4'b1001 ; B = 4'b0110 ; Cin = 1'b0 ;
#5; 
A = 4'b1001 ; B = 4'b0111 ; Cin = 1'b0 ;
#5; 
A = 4'b1001 ; B = 4'b1000 ; Cin = 1'b0 ;
#5; 
A = 4'b1001 ; B = 4'b1001 ; Cin = 1'b0 ;
#5; 
A = 4'b1001 ; B = 4'b1010 ; Cin = 1'b0 ;
#5; 
A = 4'b1001 ; B = 4'b1011 ; Cin = 1'b0 ;
#5; 
A = 4'b1001 ; B = 4'b1100 ; Cin = 1'b0 ;
#5; 
A = 4'b1001 ; B = 4'b1101 ; Cin = 1'b0 ;
#5; 
A = 4'b1001 ; B = 4'b1110 ; Cin = 1'b0 ;
#5; 
A = 4'b1001 ; B = 4'b1111 ; Cin = 1'b0 ;
#5; 
A = 4'b1010 ; B = 4'b0000 ; Cin = 1'b0 ;
#5; 
A = 4'b1010 ; B = 4'b0001 ; Cin = 1'b0 ;
#5; 
A = 4'b1010 ; B = 4'b0010 ; Cin = 1'b0 ;
#5; 
A = 4'b1010 ; B = 4'b0011 ; Cin = 1'b0 ;
#5; 
A = 4'b1010 ; B = 4'b0100 ; Cin = 1'b0 ;
#5; 
A = 4'b1010 ; B = 4'b0101 ; Cin = 1'b0 ;
#5; 
A = 4'b1010 ; B = 4'b0110 ; Cin = 1'b0 ;
#5; 
A = 4'b1010 ; B = 4'b0111 ; Cin = 1'b0 ;
#5; 
A = 4'b1010 ; B = 4'b1000 ; Cin = 1'b0 ;
#5; 
A = 4'b1010 ; B = 4'b1001 ; Cin = 1'b0 ;
#5; 
A = 4'b1010 ; B = 4'b1010 ; Cin = 1'b0 ;
#5; 
A = 4'b1010 ; B = 4'b1011 ; Cin = 1'b0 ;
#5; 
A = 4'b1010 ; B = 4'b1100 ; Cin = 1'b0 ;
#5; 
A = 4'b1010 ; B = 4'b1101 ; Cin = 1'b0 ;
#5; 
A = 4'b1010 ; B = 4'b1110 ; Cin = 1'b0 ;
#5; 
A = 4'b1010 ; B = 4'b1111 ; Cin = 1'b0 ;
#5; 
A = 4'b1011 ; B = 4'b0000 ; Cin = 1'b0 ;
#5; 
A = 4'b1011 ; B = 4'b0001 ; Cin = 1'b0 ;
#5; 
A = 4'b1011 ; B = 4'b0010 ; Cin = 1'b0 ;
#5; 
A = 4'b1011 ; B = 4'b0011 ; Cin = 1'b0 ;
#5; 
A = 4'b1011 ; B = 4'b0100 ; Cin = 1'b0 ;
#5; 
A = 4'b1011 ; B = 4'b0101 ; Cin = 1'b0 ;
#5; 
A = 4'b1011 ; B = 4'b0110 ; Cin = 1'b0 ;
#5; 
A = 4'b1011 ; B = 4'b0111 ; Cin = 1'b0 ;
#5; 
A = 4'b1011 ; B = 4'b1000 ; Cin = 1'b0 ;
#5; 
A = 4'b1011 ; B = 4'b1001 ; Cin = 1'b0 ;
#5; 
A = 4'b1011 ; B = 4'b1010 ; Cin = 1'b0 ;
#5; 
A = 4'b1011 ; B = 4'b1011 ; Cin = 1'b0 ;
#5; 
A = 4'b1011 ; B = 4'b1100 ; Cin = 1'b0 ;
#5; 
A = 4'b1011 ; B = 4'b1101 ; Cin = 1'b0 ;
#5; 
A = 4'b1011 ; B = 4'b1110 ; Cin = 1'b0 ;
#5; 
A = 4'b1011 ; B = 4'b1111 ; Cin = 1'b0 ;
#5; 
A = 4'b1100 ; B = 4'b0000 ; Cin = 1'b0 ;
#5; 
A = 4'b1100 ; B = 4'b0001 ; Cin = 1'b0 ;
#5; 
A = 4'b1100 ; B = 4'b0010 ; Cin = 1'b0 ;
#5; 
A = 4'b1100 ; B = 4'b0011 ; Cin = 1'b0 ;
#5; 
A = 4'b1100 ; B = 4'b0100 ; Cin = 1'b0 ;
#5; 
A = 4'b1100 ; B = 4'b0101 ; Cin = 1'b0 ;
#5; 
A = 4'b1100 ; B = 4'b0110 ; Cin = 1'b0 ;
#5; 
A = 4'b1100 ; B = 4'b0111 ; Cin = 1'b0 ;
#5; 
A = 4'b1100 ; B = 4'b1000 ; Cin = 1'b0 ;
#5; 
A = 4'b1100 ; B = 4'b1001 ; Cin = 1'b0 ;
#5; 
A = 4'b1100 ; B = 4'b1010 ; Cin = 1'b0 ;
#5; 
A = 4'b1100 ; B = 4'b1011 ; Cin = 1'b0 ;
#5; 
A = 4'b1100 ; B = 4'b1100 ; Cin = 1'b0 ;
#5; 
A = 4'b1100 ; B = 4'b1101 ; Cin = 1'b0 ;
#5; 
A = 4'b1100 ; B = 4'b1110 ; Cin = 1'b0 ;
#5; 
A = 4'b1100 ; B = 4'b1111 ; Cin = 1'b0 ;
#5; 
A = 4'b1101 ; B = 4'b0000 ; Cin = 1'b0 ;
#5; 
A = 4'b1101 ; B = 4'b0001 ; Cin = 1'b0 ;
#5; 
A = 4'b1101 ; B = 4'b0010 ; Cin = 1'b0 ;
#5; 
A = 4'b1101 ; B = 4'b0011 ; Cin = 1'b0 ;
#5; 
A = 4'b1101 ; B = 4'b0100 ; Cin = 1'b0 ;
#5; 
A = 4'b1101 ; B = 4'b0101 ; Cin = 1'b0 ;
#5; 
A = 4'b1101 ; B = 4'b0110 ; Cin = 1'b0 ;
#5; 
A = 4'b1101 ; B = 4'b0111 ; Cin = 1'b0 ;
#5; 
A = 4'b1101 ; B = 4'b1000 ; Cin = 1'b0 ;
#5; 
A = 4'b1101 ; B = 4'b1001 ; Cin = 1'b0 ;
#5; 
A = 4'b1101 ; B = 4'b1010 ; Cin = 1'b0 ;
#5; 
A = 4'b1101 ; B = 4'b1011 ; Cin = 1'b0 ;
#5; 
A = 4'b1101 ; B = 4'b1100 ; Cin = 1'b0 ;
#5; 
A = 4'b1101 ; B = 4'b1101 ; Cin = 1'b0 ;
#5; 
A = 4'b1101 ; B = 4'b1110 ; Cin = 1'b0 ;
#5; 
A = 4'b1101 ; B = 4'b1111 ; Cin = 1'b0 ;
#5; 
A = 4'b1110 ; B = 4'b0000 ; Cin = 1'b0 ;
#5; 
A = 4'b1110 ; B = 4'b0001 ; Cin = 1'b0 ;
#5; 
A = 4'b1110 ; B = 4'b0010 ; Cin = 1'b0 ;
#5; 
A = 4'b1110 ; B = 4'b0011 ; Cin = 1'b0 ;
#5; 
A = 4'b1110 ; B = 4'b0100 ; Cin = 1'b0 ;
#5; 
A = 4'b1110 ; B = 4'b0101 ; Cin = 1'b0 ;
#5; 
A = 4'b1110 ; B = 4'b0110 ; Cin = 1'b0 ;
#5; 
A = 4'b1110 ; B = 4'b0111 ; Cin = 1'b0 ;
#5; 
A = 4'b1110 ; B = 4'b1000 ; Cin = 1'b0 ;
#5; 
A = 4'b1110 ; B = 4'b1001 ; Cin = 1'b0 ;
#5; 
A = 4'b1110 ; B = 4'b1010 ; Cin = 1'b0 ;
#5; 
A = 4'b1110 ; B = 4'b1011 ; Cin = 1'b0 ;
#5; 
A = 4'b1110 ; B = 4'b1100 ; Cin = 1'b0 ;
#5; 
A = 4'b1110 ; B = 4'b1101 ; Cin = 1'b0 ;
#5; 
A = 4'b1110 ; B = 4'b1110 ; Cin = 1'b0 ;
#5; 
A = 4'b1110 ; B = 4'b1111 ; Cin = 1'b0 ;
#5; 
A = 4'b1111 ; B = 4'b0000 ; Cin = 1'b0 ;
#5; 
A = 4'b1111 ; B = 4'b0001 ; Cin = 1'b0 ;
#5; 
A = 4'b1111 ; B = 4'b0010 ; Cin = 1'b0 ;
#5; 
A = 4'b1111 ; B = 4'b0011 ; Cin = 1'b0 ;
#5; 
A = 4'b1111 ; B = 4'b0100 ; Cin = 1'b0 ;
#5; 
A = 4'b1111 ; B = 4'b0101 ; Cin = 1'b0 ;
#5; 
A = 4'b1111 ; B = 4'b0110 ; Cin = 1'b0 ;
#5; 
A = 4'b1111 ; B = 4'b0111 ; Cin = 1'b0 ;
#5; 
A = 4'b1111 ; B = 4'b1000 ; Cin = 1'b0 ;
#5; 
A = 4'b1111 ; B = 4'b1001 ; Cin = 1'b0 ;
#5; 
A = 4'b1111 ; B = 4'b1010 ; Cin = 1'b0 ;
#5; 
A = 4'b1111 ; B = 4'b1011 ; Cin = 1'b0 ;
#5; 
A = 4'b1111 ; B = 4'b1100 ; Cin = 1'b0 ;
#5; 
A = 4'b1111 ; B = 4'b1101 ; Cin = 1'b0 ;
#5; 
A = 4'b1111 ; B = 4'b1110 ; Cin = 1'b0 ;
#5; 
A = 4'b1111 ; B = 4'b1111 ; Cin = 1'b0 ;
#5;
A = 4'b1111 ; B = 4'b1111 ; Cin = 1'b0 ;

end
endmodule



