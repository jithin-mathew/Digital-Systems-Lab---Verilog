module full_adder(a,b,cin,sum,cout);
input a;
input b;
input cin;
output sum;
output cout;

assign sum = a^b^cin;
assign cout = (a & b) | (cin & (a^b)); 

endmodule

module bitadder(A,B,Cin,M,Sum,Cout);

input [3:0]A;
input [3:0]B;
input Cin;
input M;

output [3:0]Sum;
output Cout;

wire c1,c2,c3;
wire b0,b1,b2,b3;

assign b0 = B[0]^M;
full_adder f1(.a(A[0]),.b(b0),.cin(Cin),.sum(Sum[0]),.cout(c1));
assign b1 = B[1]^M;
full_adder f2(.a(A[1]),.b(b1),.cin(c1),.sum(Sum[1]),.cout(c2));
assign b2 = B[2]^M;
full_adder f3(.a(A[2]),.b(b2),.cin(c2),.sum(Sum[2]),.cout(c3));
assign b3 = B[3]^M;
full_adder f4(.a(A[3]),.b(b3),.cin(c3),.sum(Sum[3]),.cout(Cout));

endmodule

module testbench();
reg [3:0]A;
reg [3:0]B;
reg Cin;
reg M;
wire [3:0]Sum;
wire Cout;

bitadder tb(A,B,Cin,M,Sum,Cout);

initial
begin

$monitor("A = %b : B = %b : Cin = %b : M = %b : Sum = %b : Cout = %b ",A,B,Cin,M,Sum,Cout);
$dumpfile("4bitadder_sub.vcd");
$dumpvars;

A = 4'b0000 ; B = 4'b0000 ; Cin = 1'b0 ; M = 1'b0 ;
#5; 
A = 4'b0000 ; B = 4'b0001 ; Cin = 1'b0 ; M = 1'b0 ;
#5; 
A = 4'b0000 ; B = 4'b0010 ; Cin = 1'b0 ; M = 1'b0 ;
#5; 
A = 4'b0000 ; B = 4'b0011 ; Cin = 1'b0 ; M = 1'b0 ;
#5; 
A = 4'b0000 ; B = 4'b0100 ; Cin = 1'b0 ; M = 1'b0 ;
#5; 
A = 4'b0000 ; B = 4'b0101 ; Cin = 1'b0 ; M = 1'b0 ;
#5; 
A = 4'b0000 ; B = 4'b0110 ; Cin = 1'b0 ; M = 1'b0 ;
#5; 
A = 4'b0000 ; B = 4'b0111 ; Cin = 1'b0 ; M = 1'b0 ;
#5; 
A = 4'b0000 ; B = 4'b1000 ; Cin = 1'b0 ; M = 1'b0 ;
#5; 
A = 4'b0000 ; B = 4'b1001 ; Cin = 1'b0 ; M = 1'b0 ;
#5; 
A = 4'b0000 ; B = 4'b1010 ; Cin = 1'b0 ; M = 1'b0 ;
#5; 
A = 4'b0000 ; B = 4'b1011 ; Cin = 1'b0 ; M = 1'b0 ;
#5; 
A = 4'b0000 ; B = 4'b1100 ; Cin = 1'b0 ; M = 1'b0 ;
#5; 
A = 4'b0000 ; B = 4'b1101 ; Cin = 1'b0 ; M = 1'b0 ;
#5; 
A = 4'b0000 ; B = 4'b1110 ; Cin = 1'b0 ; M = 1'b0 ;
#5; 
A = 4'b0000 ; B = 4'b1111 ; Cin = 1'b0 ; M = 1'b0 ;
#5; 
A = 4'b0001 ; B = 4'b0000 ; Cin = 1'b0 ; M = 1'b0 ;
#5; 
A = 4'b0001 ; B = 4'b0001 ; Cin = 1'b0 ; M = 1'b0 ;
#5; 
A = 4'b0001 ; B = 4'b0010 ; Cin = 1'b0 ; M = 1'b0 ;
#5; 
A = 4'b0001 ; B = 4'b0011 ; Cin = 1'b0 ; M = 1'b0 ;
#5; 
A = 4'b0001 ; B = 4'b0100 ; Cin = 1'b0 ; M = 1'b0 ;
#5; 
A = 4'b0001 ; B = 4'b0101 ; Cin = 1'b0 ; M = 1'b0 ;
#5; 
A = 4'b0001 ; B = 4'b0110 ; Cin = 1'b0 ; M = 1'b0 ;
#5; 
A = 4'b0001 ; B = 4'b0111 ; Cin = 1'b0 ; M = 1'b0 ;
#5; 
A = 4'b0001 ; B = 4'b1000 ; Cin = 1'b0 ; M = 1'b0 ;
#5; 
A = 4'b0001 ; B = 4'b1001 ; Cin = 1'b0 ; M = 1'b0 ;
#5; 
A = 4'b0001 ; B = 4'b1010 ; Cin = 1'b0 ; M = 1'b0 ;
#5; 
A = 4'b0001 ; B = 4'b1011 ; Cin = 1'b0 ; M = 1'b0 ;
#5; 
A = 4'b0001 ; B = 4'b1100 ; Cin = 1'b0 ; M = 1'b0 ;
#5; 
A = 4'b0001 ; B = 4'b1101 ; Cin = 1'b0 ; M = 1'b0 ;
#5; 
A = 4'b0001 ; B = 4'b1110 ; Cin = 1'b0 ; M = 1'b0 ;
#5; 
A = 4'b0001 ; B = 4'b1111 ; Cin = 1'b0 ; M = 1'b0 ;
#5; 
A = 4'b0010 ; B = 4'b0000 ; Cin = 1'b0 ; M = 1'b0 ;
#5; 
A = 4'b0010 ; B = 4'b0001 ; Cin = 1'b0 ; M = 1'b0 ;
#5; 
A = 4'b0010 ; B = 4'b0010 ; Cin = 1'b0 ; M = 1'b0 ;
#5; 
A = 4'b0010 ; B = 4'b0011 ; Cin = 1'b0 ; M = 1'b0 ;
#5; 
A = 4'b0010 ; B = 4'b0100 ; Cin = 1'b0 ; M = 1'b0 ;
#5; 
A = 4'b0010 ; B = 4'b0101 ; Cin = 1'b0 ; M = 1'b0 ;
#5; 
A = 4'b0010 ; B = 4'b0110 ; Cin = 1'b0 ; M = 1'b0 ;
#5; 
A = 4'b0010 ; B = 4'b0111 ; Cin = 1'b0 ; M = 1'b0 ;
#5; 
A = 4'b0010 ; B = 4'b1000 ; Cin = 1'b0 ; M = 1'b0 ;
#5; 
A = 4'b0010 ; B = 4'b1001 ; Cin = 1'b0 ; M = 1'b0 ;
#5; 
A = 4'b0010 ; B = 4'b1010 ; Cin = 1'b0 ; M = 1'b0 ;
#5; 
A = 4'b0010 ; B = 4'b1011 ; Cin = 1'b0 ; M = 1'b0 ;
#5; 
A = 4'b0010 ; B = 4'b1100 ; Cin = 1'b0 ; M = 1'b0 ;
#5; 
A = 4'b0010 ; B = 4'b1101 ; Cin = 1'b0 ; M = 1'b0 ;
#5; 
A = 4'b0010 ; B = 4'b1110 ; Cin = 1'b0 ; M = 1'b0 ;
#5; 
A = 4'b0010 ; B = 4'b1111 ; Cin = 1'b0 ; M = 1'b0 ;
#5; 
A = 4'b0011 ; B = 4'b0000 ; Cin = 1'b0 ; M = 1'b0 ;
#5; 
A = 4'b0011 ; B = 4'b0001 ; Cin = 1'b0 ; M = 1'b0 ;
#5; 
A = 4'b0011 ; B = 4'b0010 ; Cin = 1'b0 ; M = 1'b0 ;
#5; 
A = 4'b0011 ; B = 4'b0011 ; Cin = 1'b0 ; M = 1'b0 ;
#5; 
A = 4'b0011 ; B = 4'b0100 ; Cin = 1'b0 ; M = 1'b0 ;
#5; 
A = 4'b0011 ; B = 4'b0101 ; Cin = 1'b0 ; M = 1'b0 ;
#5; 
A = 4'b0011 ; B = 4'b0110 ; Cin = 1'b0 ; M = 1'b0 ;
#5; 
A = 4'b0011 ; B = 4'b0111 ; Cin = 1'b0 ; M = 1'b0 ;
#5; 
A = 4'b0011 ; B = 4'b1000 ; Cin = 1'b0 ; M = 1'b0 ;
#5; 
A = 4'b0011 ; B = 4'b1001 ; Cin = 1'b0 ; M = 1'b0 ;
#5; 
A = 4'b0011 ; B = 4'b1010 ; Cin = 1'b0 ; M = 1'b0 ;
#5; 
A = 4'b0011 ; B = 4'b1011 ; Cin = 1'b0 ; M = 1'b0 ;
#5; 
A = 4'b0011 ; B = 4'b1100 ; Cin = 1'b0 ; M = 1'b0 ;
#5; 
A = 4'b0011 ; B = 4'b1101 ; Cin = 1'b0 ; M = 1'b0 ;
#5; 
A = 4'b0011 ; B = 4'b1110 ; Cin = 1'b0 ; M = 1'b0 ;
#5; 
A = 4'b0011 ; B = 4'b1111 ; Cin = 1'b0 ; M = 1'b0 ;
#5; 
A = 4'b0100 ; B = 4'b0000 ; Cin = 1'b0 ; M = 1'b0 ;
#5; 
A = 4'b0100 ; B = 4'b0001 ; Cin = 1'b0 ; M = 1'b0 ;
#5; 
A = 4'b0100 ; B = 4'b0010 ; Cin = 1'b0 ; M = 1'b0 ;
#5; 
A = 4'b0100 ; B = 4'b0011 ; Cin = 1'b0 ; M = 1'b0 ;
#5; 
A = 4'b0100 ; B = 4'b0100 ; Cin = 1'b0 ; M = 1'b0 ;
#5; 
A = 4'b0100 ; B = 4'b0101 ; Cin = 1'b0 ; M = 1'b0 ;
#5; 
A = 4'b0100 ; B = 4'b0110 ; Cin = 1'b0 ; M = 1'b0 ;
#5; 
A = 4'b0100 ; B = 4'b0111 ; Cin = 1'b0 ; M = 1'b0 ;
#5; 
A = 4'b0100 ; B = 4'b1000 ; Cin = 1'b0 ; M = 1'b0 ;
#5; 
A = 4'b0100 ; B = 4'b1001 ; Cin = 1'b0 ; M = 1'b0 ;
#5; 
A = 4'b0100 ; B = 4'b1010 ; Cin = 1'b0 ; M = 1'b0 ;
#5; 
A = 4'b0100 ; B = 4'b1011 ; Cin = 1'b0 ; M = 1'b0 ;
#5; 
A = 4'b0100 ; B = 4'b1100 ; Cin = 1'b0 ; M = 1'b0 ;
#5; 
A = 4'b0100 ; B = 4'b1101 ; Cin = 1'b0 ; M = 1'b0 ;
#5; 
A = 4'b0100 ; B = 4'b1110 ; Cin = 1'b0 ; M = 1'b0 ;
#5; 
A = 4'b0100 ; B = 4'b1111 ; Cin = 1'b0 ; M = 1'b0 ;
#5; 
A = 4'b0101 ; B = 4'b0000 ; Cin = 1'b0 ; M = 1'b0 ;
#5; 
A = 4'b0101 ; B = 4'b0001 ; Cin = 1'b0 ; M = 1'b0 ;
#5; 
A = 4'b0101 ; B = 4'b0010 ; Cin = 1'b0 ; M = 1'b0 ;
#5; 
A = 4'b0101 ; B = 4'b0011 ; Cin = 1'b0 ; M = 1'b0 ;
#5; 
A = 4'b0101 ; B = 4'b0100 ; Cin = 1'b0 ; M = 1'b0 ;
#5; 
A = 4'b0101 ; B = 4'b0101 ; Cin = 1'b0 ; M = 1'b0 ;
#5; 
A = 4'b0101 ; B = 4'b0110 ; Cin = 1'b0 ; M = 1'b0 ;
#5; 
A = 4'b0101 ; B = 4'b0111 ; Cin = 1'b0 ; M = 1'b0 ;
#5; 
A = 4'b0101 ; B = 4'b1000 ; Cin = 1'b0 ; M = 1'b0 ;
#5; 
A = 4'b0101 ; B = 4'b1001 ; Cin = 1'b0 ; M = 1'b0 ;
#5; 
A = 4'b0101 ; B = 4'b1010 ; Cin = 1'b0 ; M = 1'b0 ;
#5; 
A = 4'b0101 ; B = 4'b1011 ; Cin = 1'b0 ; M = 1'b0 ;
#5; 
A = 4'b0101 ; B = 4'b1100 ; Cin = 1'b0 ; M = 1'b0 ;
#5; 
A = 4'b0101 ; B = 4'b1101 ; Cin = 1'b0 ; M = 1'b0 ;
#5; 
A = 4'b0101 ; B = 4'b1110 ; Cin = 1'b0 ; M = 1'b0 ;
#5; 
A = 4'b0101 ; B = 4'b1111 ; Cin = 1'b0 ; M = 1'b0 ;
#5; 
A = 4'b0110 ; B = 4'b0000 ; Cin = 1'b0 ; M = 1'b0 ;
#5; 
A = 4'b0110 ; B = 4'b0001 ; Cin = 1'b0 ; M = 1'b0 ;
#5; 
A = 4'b0110 ; B = 4'b0010 ; Cin = 1'b0 ; M = 1'b0 ;
#5; 
A = 4'b0110 ; B = 4'b0011 ; Cin = 1'b0 ; M = 1'b0 ;
#5; 
A = 4'b0110 ; B = 4'b0100 ; Cin = 1'b0 ; M = 1'b0 ;
#5; 
A = 4'b0110 ; B = 4'b0101 ; Cin = 1'b0 ; M = 1'b0 ;
#5; 
A = 4'b0110 ; B = 4'b0110 ; Cin = 1'b0 ; M = 1'b0 ;
#5; 
A = 4'b0110 ; B = 4'b0111 ; Cin = 1'b0 ; M = 1'b0 ;
#5; 
A = 4'b0110 ; B = 4'b1000 ; Cin = 1'b0 ; M = 1'b0 ;
#5; 
A = 4'b0110 ; B = 4'b1001 ; Cin = 1'b0 ; M = 1'b0 ;
#5; 
A = 4'b0110 ; B = 4'b1010 ; Cin = 1'b0 ; M = 1'b0 ;
#5; 
A = 4'b0110 ; B = 4'b1011 ; Cin = 1'b0 ; M = 1'b0 ;
#5; 
A = 4'b0110 ; B = 4'b1100 ; Cin = 1'b0 ; M = 1'b0 ;
#5; 
A = 4'b0110 ; B = 4'b1101 ; Cin = 1'b0 ; M = 1'b0 ;
#5; 
A = 4'b0110 ; B = 4'b1110 ; Cin = 1'b0 ; M = 1'b0 ;
#5; 
A = 4'b0110 ; B = 4'b1111 ; Cin = 1'b0 ; M = 1'b0 ;
#5; 
A = 4'b0111 ; B = 4'b0000 ; Cin = 1'b0 ; M = 1'b0 ;
#5; 
A = 4'b0111 ; B = 4'b0001 ; Cin = 1'b0 ; M = 1'b0 ;
#5; 
A = 4'b0111 ; B = 4'b0010 ; Cin = 1'b0 ; M = 1'b0 ;
#5; 
A = 4'b0111 ; B = 4'b0011 ; Cin = 1'b0 ; M = 1'b0 ;
#5; 
A = 4'b0111 ; B = 4'b0100 ; Cin = 1'b0 ; M = 1'b0 ;
#5; 
A = 4'b0111 ; B = 4'b0101 ; Cin = 1'b0 ; M = 1'b0 ;
#5; 
A = 4'b0111 ; B = 4'b0110 ; Cin = 1'b0 ; M = 1'b0 ;
#5; 
A = 4'b0111 ; B = 4'b0111 ; Cin = 1'b0 ; M = 1'b0 ;
#5; 
A = 4'b0111 ; B = 4'b1000 ; Cin = 1'b0 ; M = 1'b0 ;
#5; 
A = 4'b0111 ; B = 4'b1001 ; Cin = 1'b0 ; M = 1'b0 ;
#5; 
A = 4'b0111 ; B = 4'b1010 ; Cin = 1'b0 ; M = 1'b0 ;
#5; 
A = 4'b0111 ; B = 4'b1011 ; Cin = 1'b0 ; M = 1'b0 ;
#5; 
A = 4'b0111 ; B = 4'b1100 ; Cin = 1'b0 ; M = 1'b0 ;
#5; 
A = 4'b0111 ; B = 4'b1101 ; Cin = 1'b0 ; M = 1'b0 ;
#5; 
A = 4'b0111 ; B = 4'b1110 ; Cin = 1'b0 ; M = 1'b0 ;
#5; 
A = 4'b0111 ; B = 4'b1111 ; Cin = 1'b0 ; M = 1'b0 ;
#5; 
A = 4'b1000 ; B = 4'b0000 ; Cin = 1'b0 ; M = 1'b0 ;
#5; 
A = 4'b1000 ; B = 4'b0001 ; Cin = 1'b0 ; M = 1'b0 ;
#5; 
A = 4'b1000 ; B = 4'b0010 ; Cin = 1'b0 ; M = 1'b0 ;
#5; 
A = 4'b1000 ; B = 4'b0011 ; Cin = 1'b0 ; M = 1'b0 ;
#5; 
A = 4'b1000 ; B = 4'b0100 ; Cin = 1'b0 ; M = 1'b0 ;
#5; 
A = 4'b1000 ; B = 4'b0101 ; Cin = 1'b0 ; M = 1'b0 ;
#5; 
A = 4'b1000 ; B = 4'b0110 ; Cin = 1'b0 ; M = 1'b0 ;
#5; 
A = 4'b1000 ; B = 4'b0111 ; Cin = 1'b0 ; M = 1'b0 ;
#5; 
A = 4'b1000 ; B = 4'b1000 ; Cin = 1'b0 ; M = 1'b0 ;
#5; 
A = 4'b1000 ; B = 4'b1001 ; Cin = 1'b0 ; M = 1'b0 ;
#5; 
A = 4'b1000 ; B = 4'b1010 ; Cin = 1'b0 ; M = 1'b0 ;
#5; 
A = 4'b1000 ; B = 4'b1011 ; Cin = 1'b0 ; M = 1'b0 ;
#5; 
A = 4'b1000 ; B = 4'b1100 ; Cin = 1'b0 ; M = 1'b0 ;
#5; 
A = 4'b1000 ; B = 4'b1101 ; Cin = 1'b0 ; M = 1'b0 ;
#5; 
A = 4'b1000 ; B = 4'b1110 ; Cin = 1'b0 ; M = 1'b0 ;
#5; 
A = 4'b1000 ; B = 4'b1111 ; Cin = 1'b0 ; M = 1'b0 ;
#5; 
A = 4'b1001 ; B = 4'b0000 ; Cin = 1'b0 ; M = 1'b0 ;
#5; 
A = 4'b1001 ; B = 4'b0001 ; Cin = 1'b0 ; M = 1'b0 ;
#5; 
A = 4'b1001 ; B = 4'b0010 ; Cin = 1'b0 ; M = 1'b0 ;
#5; 
A = 4'b1001 ; B = 4'b0011 ; Cin = 1'b0 ; M = 1'b0 ;
#5; 
A = 4'b1001 ; B = 4'b0100 ; Cin = 1'b0 ; M = 1'b0 ;
#5; 
A = 4'b1001 ; B = 4'b0101 ; Cin = 1'b0 ; M = 1'b0 ;
#5; 
A = 4'b1001 ; B = 4'b0110 ; Cin = 1'b0 ; M = 1'b0 ;
#5; 
A = 4'b1001 ; B = 4'b0111 ; Cin = 1'b0 ; M = 1'b0 ;
#5; 
A = 4'b1001 ; B = 4'b1000 ; Cin = 1'b0 ; M = 1'b0 ;
#5; 
A = 4'b1001 ; B = 4'b1001 ; Cin = 1'b0 ; M = 1'b0 ;
#5; 
A = 4'b1001 ; B = 4'b1010 ; Cin = 1'b0 ; M = 1'b0 ;
#5; 
A = 4'b1001 ; B = 4'b1011 ; Cin = 1'b0 ; M = 1'b0 ;
#5; 
A = 4'b1001 ; B = 4'b1100 ; Cin = 1'b0 ; M = 1'b0 ;
#5; 
A = 4'b1001 ; B = 4'b1101 ; Cin = 1'b0 ; M = 1'b0 ;
#5; 
A = 4'b1001 ; B = 4'b1110 ; Cin = 1'b0 ; M = 1'b0 ;
#5; 
A = 4'b1001 ; B = 4'b1111 ; Cin = 1'b0 ; M = 1'b0 ;
#5; 
A = 4'b1010 ; B = 4'b0000 ; Cin = 1'b0 ; M = 1'b0 ;
#5; 
A = 4'b1010 ; B = 4'b0001 ; Cin = 1'b0 ; M = 1'b0 ;
#5; 
A = 4'b1010 ; B = 4'b0010 ; Cin = 1'b0 ; M = 1'b0 ;
#5; 
A = 4'b1010 ; B = 4'b0011 ; Cin = 1'b0 ; M = 1'b0 ;
#5; 
A = 4'b1010 ; B = 4'b0100 ; Cin = 1'b0 ; M = 1'b0 ;
#5; 
A = 4'b1010 ; B = 4'b0101 ; Cin = 1'b0 ; M = 1'b0 ;
#5; 
A = 4'b1010 ; B = 4'b0110 ; Cin = 1'b0 ; M = 1'b0 ;
#5; 
A = 4'b1010 ; B = 4'b0111 ; Cin = 1'b0 ; M = 1'b0 ;
#5; 
A = 4'b1010 ; B = 4'b1000 ; Cin = 1'b0 ; M = 1'b0 ;
#5; 
A = 4'b1010 ; B = 4'b1001 ; Cin = 1'b0 ; M = 1'b0 ;
#5; 
A = 4'b1010 ; B = 4'b1010 ; Cin = 1'b0 ; M = 1'b0 ;
#5; 
A = 4'b1010 ; B = 4'b1011 ; Cin = 1'b0 ; M = 1'b0 ;
#5; 
A = 4'b1010 ; B = 4'b1100 ; Cin = 1'b0 ; M = 1'b0 ;
#5; 
A = 4'b1010 ; B = 4'b1101 ; Cin = 1'b0 ; M = 1'b0 ;
#5; 
A = 4'b1010 ; B = 4'b1110 ; Cin = 1'b0 ; M = 1'b0 ;
#5; 
A = 4'b1010 ; B = 4'b1111 ; Cin = 1'b0 ; M = 1'b0 ;
#5; 
A = 4'b1011 ; B = 4'b0000 ; Cin = 1'b0 ; M = 1'b0 ;
#5; 
A = 4'b1011 ; B = 4'b0001 ; Cin = 1'b0 ; M = 1'b0 ;
#5; 
A = 4'b1011 ; B = 4'b0010 ; Cin = 1'b0 ; M = 1'b0 ;
#5; 
A = 4'b1011 ; B = 4'b0011 ; Cin = 1'b0 ; M = 1'b0 ;
#5; 
A = 4'b1011 ; B = 4'b0100 ; Cin = 1'b0 ; M = 1'b0 ;
#5; 
A = 4'b1011 ; B = 4'b0101 ; Cin = 1'b0 ; M = 1'b0 ;
#5; 
A = 4'b1011 ; B = 4'b0110 ; Cin = 1'b0 ; M = 1'b0 ;
#5; 
A = 4'b1011 ; B = 4'b0111 ; Cin = 1'b0 ; M = 1'b0 ;
#5; 
A = 4'b1011 ; B = 4'b1000 ; Cin = 1'b0 ; M = 1'b0 ;
#5; 
A = 4'b1011 ; B = 4'b1001 ; Cin = 1'b0 ; M = 1'b0 ;
#5; 
A = 4'b1011 ; B = 4'b1010 ; Cin = 1'b0 ; M = 1'b0 ;
#5; 
A = 4'b1011 ; B = 4'b1011 ; Cin = 1'b0 ; M = 1'b0 ;
#5; 
A = 4'b1011 ; B = 4'b1100 ; Cin = 1'b0 ; M = 1'b0 ;
#5; 
A = 4'b1011 ; B = 4'b1101 ; Cin = 1'b0 ; M = 1'b0 ;
#5; 
A = 4'b1011 ; B = 4'b1110 ; Cin = 1'b0 ; M = 1'b0 ;
#5; 
A = 4'b1011 ; B = 4'b1111 ; Cin = 1'b0 ; M = 1'b0 ;
#5; 
A = 4'b1100 ; B = 4'b0000 ; Cin = 1'b0 ; M = 1'b0 ;
#5; 
A = 4'b1100 ; B = 4'b0001 ; Cin = 1'b0 ; M = 1'b0 ;
#5; 
A = 4'b1100 ; B = 4'b0010 ; Cin = 1'b0 ; M = 1'b0 ;
#5; 
A = 4'b1100 ; B = 4'b0011 ; Cin = 1'b0 ; M = 1'b0 ;
#5; 
A = 4'b1100 ; B = 4'b0100 ; Cin = 1'b0 ; M = 1'b0 ;
#5; 
A = 4'b1100 ; B = 4'b0101 ; Cin = 1'b0 ; M = 1'b0 ;
#5; 
A = 4'b1100 ; B = 4'b0110 ; Cin = 1'b0 ; M = 1'b0 ;
#5; 
A = 4'b1100 ; B = 4'b0111 ; Cin = 1'b0 ; M = 1'b0 ;
#5; 
A = 4'b1100 ; B = 4'b1000 ; Cin = 1'b0 ; M = 1'b0 ;
#5; 
A = 4'b1100 ; B = 4'b1001 ; Cin = 1'b0 ; M = 1'b0 ;
#5; 
A = 4'b1100 ; B = 4'b1010 ; Cin = 1'b0 ; M = 1'b0 ;
#5; 
A = 4'b1100 ; B = 4'b1011 ; Cin = 1'b0 ; M = 1'b0 ;
#5; 
A = 4'b1100 ; B = 4'b1100 ; Cin = 1'b0 ; M = 1'b0 ;
#5; 
A = 4'b1100 ; B = 4'b1101 ; Cin = 1'b0 ; M = 1'b0 ;
#5; 
A = 4'b1100 ; B = 4'b1110 ; Cin = 1'b0 ; M = 1'b0 ;
#5; 
A = 4'b1100 ; B = 4'b1111 ; Cin = 1'b0 ; M = 1'b0 ;
#5; 
A = 4'b1101 ; B = 4'b0000 ; Cin = 1'b0 ; M = 1'b0 ;
#5; 
A = 4'b1101 ; B = 4'b0001 ; Cin = 1'b0 ; M = 1'b0 ;
#5; 
A = 4'b1101 ; B = 4'b0010 ; Cin = 1'b0 ; M = 1'b0 ;
#5; 
A = 4'b1101 ; B = 4'b0011 ; Cin = 1'b0 ; M = 1'b0 ;
#5; 
A = 4'b1101 ; B = 4'b0100 ; Cin = 1'b0 ; M = 1'b0 ;
#5; 
A = 4'b1101 ; B = 4'b0101 ; Cin = 1'b0 ; M = 1'b0 ;
#5; 
A = 4'b1101 ; B = 4'b0110 ; Cin = 1'b0 ; M = 1'b0 ;
#5; 
A = 4'b1101 ; B = 4'b0111 ; Cin = 1'b0 ; M = 1'b0 ;
#5; 
A = 4'b1101 ; B = 4'b1000 ; Cin = 1'b0 ; M = 1'b0 ;
#5; 
A = 4'b1101 ; B = 4'b1001 ; Cin = 1'b0 ; M = 1'b0 ;
#5; 
A = 4'b1101 ; B = 4'b1010 ; Cin = 1'b0 ; M = 1'b0 ;
#5; 
A = 4'b1101 ; B = 4'b1011 ; Cin = 1'b0 ; M = 1'b0 ;
#5; 
A = 4'b1101 ; B = 4'b1100 ; Cin = 1'b0 ; M = 1'b0 ;
#5; 
A = 4'b1101 ; B = 4'b1101 ; Cin = 1'b0 ; M = 1'b0 ;
#5; 
A = 4'b1101 ; B = 4'b1110 ; Cin = 1'b0 ; M = 1'b0 ;
#5; 
A = 4'b1101 ; B = 4'b1111 ; Cin = 1'b0 ; M = 1'b0 ;
#5; 
A = 4'b1110 ; B = 4'b0000 ; Cin = 1'b0 ; M = 1'b0 ;
#5; 
A = 4'b1110 ; B = 4'b0001 ; Cin = 1'b0 ; M = 1'b0 ;
#5; 
A = 4'b1110 ; B = 4'b0010 ; Cin = 1'b0 ; M = 1'b0 ;
#5; 
A = 4'b1110 ; B = 4'b0011 ; Cin = 1'b0 ; M = 1'b0 ;
#5; 
A = 4'b1110 ; B = 4'b0100 ; Cin = 1'b0 ; M = 1'b0 ;
#5; 
A = 4'b1110 ; B = 4'b0101 ; Cin = 1'b0 ; M = 1'b0 ;
#5; 
A = 4'b1110 ; B = 4'b0110 ; Cin = 1'b0 ; M = 1'b0 ;
#5; 
A = 4'b1110 ; B = 4'b0111 ; Cin = 1'b0 ; M = 1'b0 ;
#5; 
A = 4'b1110 ; B = 4'b1000 ; Cin = 1'b0 ; M = 1'b0 ;
#5; 
A = 4'b1110 ; B = 4'b1001 ; Cin = 1'b0 ; M = 1'b0 ;
#5; 
A = 4'b1110 ; B = 4'b1010 ; Cin = 1'b0 ; M = 1'b0 ;
#5; 
A = 4'b1110 ; B = 4'b1011 ; Cin = 1'b0 ; M = 1'b0 ;
#5; 
A = 4'b1110 ; B = 4'b1100 ; Cin = 1'b0 ; M = 1'b0 ;
#5; 
A = 4'b1110 ; B = 4'b1101 ; Cin = 1'b0 ; M = 1'b0 ;
#5; 
A = 4'b1110 ; B = 4'b1110 ; Cin = 1'b0 ; M = 1'b0 ;
#5; 
A = 4'b1110 ; B = 4'b1111 ; Cin = 1'b0 ; M = 1'b0 ;
#5; 
A = 4'b1111 ; B = 4'b0000 ; Cin = 1'b0 ; M = 1'b0 ;
#5; 
A = 4'b1111 ; B = 4'b0001 ; Cin = 1'b0 ; M = 1'b0 ;
#5; 
A = 4'b1111 ; B = 4'b0010 ; Cin = 1'b0 ; M = 1'b0 ;
#5; 
A = 4'b1111 ; B = 4'b0011 ; Cin = 1'b0 ; M = 1'b0 ;
#5; 
A = 4'b1111 ; B = 4'b0100 ; Cin = 1'b0 ; M = 1'b0 ;
#5; 
A = 4'b1111 ; B = 4'b0101 ; Cin = 1'b0 ; M = 1'b0 ;
#5; 
A = 4'b1111 ; B = 4'b0110 ; Cin = 1'b0 ; M = 1'b0 ;
#5; 
A = 4'b1111 ; B = 4'b0111 ; Cin = 1'b0 ; M = 1'b0 ;
#5; 
A = 4'b1111 ; B = 4'b1000 ; Cin = 1'b0 ; M = 1'b0 ;
#5; 
A = 4'b1111 ; B = 4'b1001 ; Cin = 1'b0 ; M = 1'b0 ;
#5; 
A = 4'b1111 ; B = 4'b1010 ; Cin = 1'b0 ; M = 1'b0 ;
#5; 
A = 4'b1111 ; B = 4'b1011 ; Cin = 1'b0 ; M = 1'b0 ;
#5; 
A = 4'b1111 ; B = 4'b1100 ; Cin = 1'b0 ; M = 1'b0 ;
#5; 
A = 4'b1111 ; B = 4'b1101 ; Cin = 1'b0 ; M = 1'b0 ;
#5; 
A = 4'b1111 ; B = 4'b1110 ; Cin = 1'b0 ; M = 1'b0 ;
#5; 
A = 4'b1111 ; B = 4'b1111 ; Cin = 1'b0 ; M = 1'b0 ;
#5; 
A = 4'b0000 ; B = 4'b0000 ; Cin = 1'b0 ; M = 1'b1 ;
#5; 
A = 4'b0000 ; B = 4'b0001 ; Cin = 1'b0 ; M = 1'b1 ;
#5; 
A = 4'b0000 ; B = 4'b0010 ; Cin = 1'b0 ; M = 1'b1 ;
#5; 
A = 4'b0000 ; B = 4'b0011 ; Cin = 1'b0 ; M = 1'b1 ;
#5; 
A = 4'b0000 ; B = 4'b0100 ; Cin = 1'b0 ; M = 1'b1 ;
#5; 
A = 4'b0000 ; B = 4'b0101 ; Cin = 1'b0 ; M = 1'b1 ;
#5; 
A = 4'b0000 ; B = 4'b0110 ; Cin = 1'b0 ; M = 1'b1 ;
#5; 
A = 4'b0000 ; B = 4'b0111 ; Cin = 1'b0 ; M = 1'b1 ;
#5; 
A = 4'b0000 ; B = 4'b1000 ; Cin = 1'b0 ; M = 1'b1 ;
#5; 
A = 4'b0000 ; B = 4'b1001 ; Cin = 1'b0 ; M = 1'b1 ;
#5; 
A = 4'b0000 ; B = 4'b1010 ; Cin = 1'b0 ; M = 1'b1 ;
#5; 
A = 4'b0000 ; B = 4'b1011 ; Cin = 1'b0 ; M = 1'b1 ;
#5; 
A = 4'b0000 ; B = 4'b1100 ; Cin = 1'b0 ; M = 1'b1 ;
#5; 
A = 4'b0000 ; B = 4'b1101 ; Cin = 1'b0 ; M = 1'b1 ;
#5; 
A = 4'b0000 ; B = 4'b1110 ; Cin = 1'b0 ; M = 1'b1 ;
#5; 
A = 4'b0000 ; B = 4'b1111 ; Cin = 1'b0 ; M = 1'b1 ;
#5; 
A = 4'b0001 ; B = 4'b0000 ; Cin = 1'b0 ; M = 1'b1 ;
#5; 
A = 4'b0001 ; B = 4'b0001 ; Cin = 1'b0 ; M = 1'b1 ;
#5; 
A = 4'b0001 ; B = 4'b0010 ; Cin = 1'b0 ; M = 1'b1 ;
#5; 
A = 4'b0001 ; B = 4'b0011 ; Cin = 1'b0 ; M = 1'b1 ;
#5; 
A = 4'b0001 ; B = 4'b0100 ; Cin = 1'b0 ; M = 1'b1 ;
#5; 
A = 4'b0001 ; B = 4'b0101 ; Cin = 1'b0 ; M = 1'b1 ;
#5; 
A = 4'b0001 ; B = 4'b0110 ; Cin = 1'b0 ; M = 1'b1 ;
#5; 
A = 4'b0001 ; B = 4'b0111 ; Cin = 1'b0 ; M = 1'b1 ;
#5; 
A = 4'b0001 ; B = 4'b1000 ; Cin = 1'b0 ; M = 1'b1 ;
#5; 
A = 4'b0001 ; B = 4'b1001 ; Cin = 1'b0 ; M = 1'b1 ;
#5; 
A = 4'b0001 ; B = 4'b1010 ; Cin = 1'b0 ; M = 1'b1 ;
#5; 
A = 4'b0001 ; B = 4'b1011 ; Cin = 1'b0 ; M = 1'b1 ;
#5; 
A = 4'b0001 ; B = 4'b1100 ; Cin = 1'b0 ; M = 1'b1 ;
#5; 
A = 4'b0001 ; B = 4'b1101 ; Cin = 1'b0 ; M = 1'b1 ;
#5; 
A = 4'b0001 ; B = 4'b1110 ; Cin = 1'b0 ; M = 1'b1 ;
#5; 
A = 4'b0001 ; B = 4'b1111 ; Cin = 1'b0 ; M = 1'b1 ;
#5; 
A = 4'b0010 ; B = 4'b0000 ; Cin = 1'b0 ; M = 1'b1 ;
#5; 
A = 4'b0010 ; B = 4'b0001 ; Cin = 1'b0 ; M = 1'b1 ;
#5; 
A = 4'b0010 ; B = 4'b0010 ; Cin = 1'b0 ; M = 1'b1 ;
#5; 
A = 4'b0010 ; B = 4'b0011 ; Cin = 1'b0 ; M = 1'b1 ;
#5; 
A = 4'b0010 ; B = 4'b0100 ; Cin = 1'b0 ; M = 1'b1 ;
#5; 
A = 4'b0010 ; B = 4'b0101 ; Cin = 1'b0 ; M = 1'b1 ;
#5; 
A = 4'b0010 ; B = 4'b0110 ; Cin = 1'b0 ; M = 1'b1 ;
#5; 
A = 4'b0010 ; B = 4'b0111 ; Cin = 1'b0 ; M = 1'b1 ;
#5; 
A = 4'b0010 ; B = 4'b1000 ; Cin = 1'b0 ; M = 1'b1 ;
#5; 
A = 4'b0010 ; B = 4'b1001 ; Cin = 1'b0 ; M = 1'b1 ;
#5; 
A = 4'b0010 ; B = 4'b1010 ; Cin = 1'b0 ; M = 1'b1 ;
#5; 
A = 4'b0010 ; B = 4'b1011 ; Cin = 1'b0 ; M = 1'b1 ;
#5; 
A = 4'b0010 ; B = 4'b1100 ; Cin = 1'b0 ; M = 1'b1 ;
#5; 
A = 4'b0010 ; B = 4'b1101 ; Cin = 1'b0 ; M = 1'b1 ;
#5; 
A = 4'b0010 ; B = 4'b1110 ; Cin = 1'b0 ; M = 1'b1 ;
#5; 
A = 4'b0010 ; B = 4'b1111 ; Cin = 1'b0 ; M = 1'b1 ;
#5; 
A = 4'b0011 ; B = 4'b0000 ; Cin = 1'b0 ; M = 1'b1 ;
#5; 
A = 4'b0011 ; B = 4'b0001 ; Cin = 1'b0 ; M = 1'b1 ;
#5; 
A = 4'b0011 ; B = 4'b0010 ; Cin = 1'b0 ; M = 1'b1 ;
#5; 
A = 4'b0011 ; B = 4'b0011 ; Cin = 1'b0 ; M = 1'b1 ;
#5; 
A = 4'b0011 ; B = 4'b0100 ; Cin = 1'b0 ; M = 1'b1 ;
#5; 
A = 4'b0011 ; B = 4'b0101 ; Cin = 1'b0 ; M = 1'b1 ;
#5; 
A = 4'b0011 ; B = 4'b0110 ; Cin = 1'b0 ; M = 1'b1 ;
#5; 
A = 4'b0011 ; B = 4'b0111 ; Cin = 1'b0 ; M = 1'b1 ;
#5; 
A = 4'b0011 ; B = 4'b1000 ; Cin = 1'b0 ; M = 1'b1 ;
#5; 
A = 4'b0011 ; B = 4'b1001 ; Cin = 1'b0 ; M = 1'b1 ;
#5; 
A = 4'b0011 ; B = 4'b1010 ; Cin = 1'b0 ; M = 1'b1 ;
#5; 
A = 4'b0011 ; B = 4'b1011 ; Cin = 1'b0 ; M = 1'b1 ;
#5; 
A = 4'b0011 ; B = 4'b1100 ; Cin = 1'b0 ; M = 1'b1 ;
#5; 
A = 4'b0011 ; B = 4'b1101 ; Cin = 1'b0 ; M = 1'b1 ;
#5; 
A = 4'b0011 ; B = 4'b1110 ; Cin = 1'b0 ; M = 1'b1 ;
#5; 
A = 4'b0011 ; B = 4'b1111 ; Cin = 1'b0 ; M = 1'b1 ;
#5; 
A = 4'b0100 ; B = 4'b0000 ; Cin = 1'b0 ; M = 1'b1 ;
#5; 
A = 4'b0100 ; B = 4'b0001 ; Cin = 1'b0 ; M = 1'b1 ;
#5; 
A = 4'b0100 ; B = 4'b0010 ; Cin = 1'b0 ; M = 1'b1 ;
#5; 
A = 4'b0100 ; B = 4'b0011 ; Cin = 1'b0 ; M = 1'b1 ;
#5; 
A = 4'b0100 ; B = 4'b0100 ; Cin = 1'b0 ; M = 1'b1 ;
#5; 
A = 4'b0100 ; B = 4'b0101 ; Cin = 1'b0 ; M = 1'b1 ;
#5; 
A = 4'b0100 ; B = 4'b0110 ; Cin = 1'b0 ; M = 1'b1 ;
#5; 
A = 4'b0100 ; B = 4'b0111 ; Cin = 1'b0 ; M = 1'b1 ;
#5; 
A = 4'b0100 ; B = 4'b1000 ; Cin = 1'b0 ; M = 1'b1 ;
#5; 
A = 4'b0100 ; B = 4'b1001 ; Cin = 1'b0 ; M = 1'b1 ;
#5; 
A = 4'b0100 ; B = 4'b1010 ; Cin = 1'b0 ; M = 1'b1 ;
#5; 
A = 4'b0100 ; B = 4'b1011 ; Cin = 1'b0 ; M = 1'b1 ;
#5; 
A = 4'b0100 ; B = 4'b1100 ; Cin = 1'b0 ; M = 1'b1 ;
#5; 
A = 4'b0100 ; B = 4'b1101 ; Cin = 1'b0 ; M = 1'b1 ;
#5; 
A = 4'b0100 ; B = 4'b1110 ; Cin = 1'b0 ; M = 1'b1 ;
#5; 
A = 4'b0100 ; B = 4'b1111 ; Cin = 1'b0 ; M = 1'b1 ;
#5; 
A = 4'b0101 ; B = 4'b0000 ; Cin = 1'b0 ; M = 1'b1 ;
#5; 
A = 4'b0101 ; B = 4'b0001 ; Cin = 1'b0 ; M = 1'b1 ;
#5; 
A = 4'b0101 ; B = 4'b0010 ; Cin = 1'b0 ; M = 1'b1 ;
#5; 
A = 4'b0101 ; B = 4'b0011 ; Cin = 1'b0 ; M = 1'b1 ;
#5; 
A = 4'b0101 ; B = 4'b0100 ; Cin = 1'b0 ; M = 1'b1 ;
#5; 
A = 4'b0101 ; B = 4'b0101 ; Cin = 1'b0 ; M = 1'b1 ;
#5; 
A = 4'b0101 ; B = 4'b0110 ; Cin = 1'b0 ; M = 1'b1 ;
#5; 
A = 4'b0101 ; B = 4'b0111 ; Cin = 1'b0 ; M = 1'b1 ;
#5; 
A = 4'b0101 ; B = 4'b1000 ; Cin = 1'b0 ; M = 1'b1 ;
#5; 
A = 4'b0101 ; B = 4'b1001 ; Cin = 1'b0 ; M = 1'b1 ;
#5; 
A = 4'b0101 ; B = 4'b1010 ; Cin = 1'b0 ; M = 1'b1 ;
#5; 
A = 4'b0101 ; B = 4'b1011 ; Cin = 1'b0 ; M = 1'b1 ;
#5; 
A = 4'b0101 ; B = 4'b1100 ; Cin = 1'b0 ; M = 1'b1 ;
#5; 
A = 4'b0101 ; B = 4'b1101 ; Cin = 1'b0 ; M = 1'b1 ;
#5; 
A = 4'b0101 ; B = 4'b1110 ; Cin = 1'b0 ; M = 1'b1 ;
#5; 
A = 4'b0101 ; B = 4'b1111 ; Cin = 1'b0 ; M = 1'b1 ;
#5; 
A = 4'b0110 ; B = 4'b0000 ; Cin = 1'b0 ; M = 1'b1 ;
#5; 
A = 4'b0110 ; B = 4'b0001 ; Cin = 1'b0 ; M = 1'b1 ;
#5; 
A = 4'b0110 ; B = 4'b0010 ; Cin = 1'b0 ; M = 1'b1 ;
#5; 
A = 4'b0110 ; B = 4'b0011 ; Cin = 1'b0 ; M = 1'b1 ;
#5; 
A = 4'b0110 ; B = 4'b0100 ; Cin = 1'b0 ; M = 1'b1 ;
#5; 
A = 4'b0110 ; B = 4'b0101 ; Cin = 1'b0 ; M = 1'b1 ;
#5; 
A = 4'b0110 ; B = 4'b0110 ; Cin = 1'b0 ; M = 1'b1 ;
#5; 
A = 4'b0110 ; B = 4'b0111 ; Cin = 1'b0 ; M = 1'b1 ;
#5; 
A = 4'b0110 ; B = 4'b1000 ; Cin = 1'b0 ; M = 1'b1 ;
#5; 
A = 4'b0110 ; B = 4'b1001 ; Cin = 1'b0 ; M = 1'b1 ;
#5; 
A = 4'b0110 ; B = 4'b1010 ; Cin = 1'b0 ; M = 1'b1 ;
#5; 
A = 4'b0110 ; B = 4'b1011 ; Cin = 1'b0 ; M = 1'b1 ;
#5; 
A = 4'b0110 ; B = 4'b1100 ; Cin = 1'b0 ; M = 1'b1 ;
#5; 
A = 4'b0110 ; B = 4'b1101 ; Cin = 1'b0 ; M = 1'b1 ;
#5; 
A = 4'b0110 ; B = 4'b1110 ; Cin = 1'b0 ; M = 1'b1 ;
#5; 
A = 4'b0110 ; B = 4'b1111 ; Cin = 1'b0 ; M = 1'b1 ;
#5; 
A = 4'b0111 ; B = 4'b0000 ; Cin = 1'b0 ; M = 1'b1 ;
#5; 
A = 4'b0111 ; B = 4'b0001 ; Cin = 1'b0 ; M = 1'b1 ;
#5; 
A = 4'b0111 ; B = 4'b0010 ; Cin = 1'b0 ; M = 1'b1 ;
#5; 
A = 4'b0111 ; B = 4'b0011 ; Cin = 1'b0 ; M = 1'b1 ;
#5; 
A = 4'b0111 ; B = 4'b0100 ; Cin = 1'b0 ; M = 1'b1 ;
#5; 
A = 4'b0111 ; B = 4'b0101 ; Cin = 1'b0 ; M = 1'b1 ;
#5; 
A = 4'b0111 ; B = 4'b0110 ; Cin = 1'b0 ; M = 1'b1 ;
#5; 
A = 4'b0111 ; B = 4'b0111 ; Cin = 1'b0 ; M = 1'b1 ;
#5; 
A = 4'b0111 ; B = 4'b1000 ; Cin = 1'b0 ; M = 1'b1 ;
#5; 
A = 4'b0111 ; B = 4'b1001 ; Cin = 1'b0 ; M = 1'b1 ;
#5; 
A = 4'b0111 ; B = 4'b1010 ; Cin = 1'b0 ; M = 1'b1 ;
#5; 
A = 4'b0111 ; B = 4'b1011 ; Cin = 1'b0 ; M = 1'b1 ;
#5; 
A = 4'b0111 ; B = 4'b1100 ; Cin = 1'b0 ; M = 1'b1 ;
#5; 
A = 4'b0111 ; B = 4'b1101 ; Cin = 1'b0 ; M = 1'b1 ;
#5; 
A = 4'b0111 ; B = 4'b1110 ; Cin = 1'b0 ; M = 1'b1 ;
#5; 
A = 4'b0111 ; B = 4'b1111 ; Cin = 1'b0 ; M = 1'b1 ;
#5; 
A = 4'b1000 ; B = 4'b0000 ; Cin = 1'b0 ; M = 1'b1 ;
#5; 
A = 4'b1000 ; B = 4'b0001 ; Cin = 1'b0 ; M = 1'b1 ;
#5; 
A = 4'b1000 ; B = 4'b0010 ; Cin = 1'b0 ; M = 1'b1 ;
#5; 
A = 4'b1000 ; B = 4'b0011 ; Cin = 1'b0 ; M = 1'b1 ;
#5; 
A = 4'b1000 ; B = 4'b0100 ; Cin = 1'b0 ; M = 1'b1 ;
#5; 
A = 4'b1000 ; B = 4'b0101 ; Cin = 1'b0 ; M = 1'b1 ;
#5; 
A = 4'b1000 ; B = 4'b0110 ; Cin = 1'b0 ; M = 1'b1 ;
#5; 
A = 4'b1000 ; B = 4'b0111 ; Cin = 1'b0 ; M = 1'b1 ;
#5; 
A = 4'b1000 ; B = 4'b1000 ; Cin = 1'b0 ; M = 1'b1 ;
#5; 
A = 4'b1000 ; B = 4'b1001 ; Cin = 1'b0 ; M = 1'b1 ;
#5; 
A = 4'b1000 ; B = 4'b1010 ; Cin = 1'b0 ; M = 1'b1 ;
#5; 
A = 4'b1000 ; B = 4'b1011 ; Cin = 1'b0 ; M = 1'b1 ;
#5; 
A = 4'b1000 ; B = 4'b1100 ; Cin = 1'b0 ; M = 1'b1 ;
#5; 
A = 4'b1000 ; B = 4'b1101 ; Cin = 1'b0 ; M = 1'b1 ;
#5; 
A = 4'b1000 ; B = 4'b1110 ; Cin = 1'b0 ; M = 1'b1 ;
#5; 
A = 4'b1000 ; B = 4'b1111 ; Cin = 1'b0 ; M = 1'b1 ;
#5; 
A = 4'b1001 ; B = 4'b0000 ; Cin = 1'b0 ; M = 1'b1 ;
#5; 
A = 4'b1001 ; B = 4'b0001 ; Cin = 1'b0 ; M = 1'b1 ;
#5; 
A = 4'b1001 ; B = 4'b0010 ; Cin = 1'b0 ; M = 1'b1 ;
#5; 
A = 4'b1001 ; B = 4'b0011 ; Cin = 1'b0 ; M = 1'b1 ;
#5; 
A = 4'b1001 ; B = 4'b0100 ; Cin = 1'b0 ; M = 1'b1 ;
#5; 
A = 4'b1001 ; B = 4'b0101 ; Cin = 1'b0 ; M = 1'b1 ;
#5; 
A = 4'b1001 ; B = 4'b0110 ; Cin = 1'b0 ; M = 1'b1 ;
#5; 
A = 4'b1001 ; B = 4'b0111 ; Cin = 1'b0 ; M = 1'b1 ;
#5; 
A = 4'b1001 ; B = 4'b1000 ; Cin = 1'b0 ; M = 1'b1 ;
#5; 
A = 4'b1001 ; B = 4'b1001 ; Cin = 1'b0 ; M = 1'b1 ;
#5; 
A = 4'b1001 ; B = 4'b1010 ; Cin = 1'b0 ; M = 1'b1 ;
#5; 
A = 4'b1001 ; B = 4'b1011 ; Cin = 1'b0 ; M = 1'b1 ;
#5; 
A = 4'b1001 ; B = 4'b1100 ; Cin = 1'b0 ; M = 1'b1 ;
#5; 
A = 4'b1001 ; B = 4'b1101 ; Cin = 1'b0 ; M = 1'b1 ;
#5; 
A = 4'b1001 ; B = 4'b1110 ; Cin = 1'b0 ; M = 1'b1 ;
#5; 
A = 4'b1001 ; B = 4'b1111 ; Cin = 1'b0 ; M = 1'b1 ;
#5; 
A = 4'b1010 ; B = 4'b0000 ; Cin = 1'b0 ; M = 1'b1 ;
#5; 
A = 4'b1010 ; B = 4'b0001 ; Cin = 1'b0 ; M = 1'b1 ;
#5; 
A = 4'b1010 ; B = 4'b0010 ; Cin = 1'b0 ; M = 1'b1 ;
#5; 
A = 4'b1010 ; B = 4'b0011 ; Cin = 1'b0 ; M = 1'b1 ;
#5; 
A = 4'b1010 ; B = 4'b0100 ; Cin = 1'b0 ; M = 1'b1 ;
#5; 
A = 4'b1010 ; B = 4'b0101 ; Cin = 1'b0 ; M = 1'b1 ;
#5; 
A = 4'b1010 ; B = 4'b0110 ; Cin = 1'b0 ; M = 1'b1 ;
#5; 
A = 4'b1010 ; B = 4'b0111 ; Cin = 1'b0 ; M = 1'b1 ;
#5; 
A = 4'b1010 ; B = 4'b1000 ; Cin = 1'b0 ; M = 1'b1 ;
#5; 
A = 4'b1010 ; B = 4'b1001 ; Cin = 1'b0 ; M = 1'b1 ;
#5; 
A = 4'b1010 ; B = 4'b1010 ; Cin = 1'b0 ; M = 1'b1 ;
#5; 
A = 4'b1010 ; B = 4'b1011 ; Cin = 1'b0 ; M = 1'b1 ;
#5; 
A = 4'b1010 ; B = 4'b1100 ; Cin = 1'b0 ; M = 1'b1 ;
#5; 
A = 4'b1010 ; B = 4'b1101 ; Cin = 1'b0 ; M = 1'b1 ;
#5; 
A = 4'b1010 ; B = 4'b1110 ; Cin = 1'b0 ; M = 1'b1 ;
#5; 
A = 4'b1010 ; B = 4'b1111 ; Cin = 1'b0 ; M = 1'b1 ;
#5; 
A = 4'b1011 ; B = 4'b0000 ; Cin = 1'b0 ; M = 1'b1 ;
#5; 
A = 4'b1011 ; B = 4'b0001 ; Cin = 1'b0 ; M = 1'b1 ;
#5; 
A = 4'b1011 ; B = 4'b0010 ; Cin = 1'b0 ; M = 1'b1 ;
#5; 
A = 4'b1011 ; B = 4'b0011 ; Cin = 1'b0 ; M = 1'b1 ;
#5; 
A = 4'b1011 ; B = 4'b0100 ; Cin = 1'b0 ; M = 1'b1 ;
#5; 
A = 4'b1011 ; B = 4'b0101 ; Cin = 1'b0 ; M = 1'b1 ;
#5; 
A = 4'b1011 ; B = 4'b0110 ; Cin = 1'b0 ; M = 1'b1 ;
#5; 
A = 4'b1011 ; B = 4'b0111 ; Cin = 1'b0 ; M = 1'b1 ;
#5; 
A = 4'b1011 ; B = 4'b1000 ; Cin = 1'b0 ; M = 1'b1 ;
#5; 
A = 4'b1011 ; B = 4'b1001 ; Cin = 1'b0 ; M = 1'b1 ;
#5; 
A = 4'b1011 ; B = 4'b1010 ; Cin = 1'b0 ; M = 1'b1 ;
#5; 
A = 4'b1011 ; B = 4'b1011 ; Cin = 1'b0 ; M = 1'b1 ;
#5; 
A = 4'b1011 ; B = 4'b1100 ; Cin = 1'b0 ; M = 1'b1 ;
#5; 
A = 4'b1011 ; B = 4'b1101 ; Cin = 1'b0 ; M = 1'b1 ;
#5; 
A = 4'b1011 ; B = 4'b1110 ; Cin = 1'b0 ; M = 1'b1 ;
#5; 
A = 4'b1011 ; B = 4'b1111 ; Cin = 1'b0 ; M = 1'b1 ;
#5; 
A = 4'b1100 ; B = 4'b0000 ; Cin = 1'b0 ; M = 1'b1 ;
#5; 
A = 4'b1100 ; B = 4'b0001 ; Cin = 1'b0 ; M = 1'b1 ;
#5; 
A = 4'b1100 ; B = 4'b0010 ; Cin = 1'b0 ; M = 1'b1 ;
#5; 
A = 4'b1100 ; B = 4'b0011 ; Cin = 1'b0 ; M = 1'b1 ;
#5; 
A = 4'b1100 ; B = 4'b0100 ; Cin = 1'b0 ; M = 1'b1 ;
#5; 
A = 4'b1100 ; B = 4'b0101 ; Cin = 1'b0 ; M = 1'b1 ;
#5; 
A = 4'b1100 ; B = 4'b0110 ; Cin = 1'b0 ; M = 1'b1 ;
#5; 
A = 4'b1100 ; B = 4'b0111 ; Cin = 1'b0 ; M = 1'b1 ;
#5; 
A = 4'b1100 ; B = 4'b1000 ; Cin = 1'b0 ; M = 1'b1 ;
#5; 
A = 4'b1100 ; B = 4'b1001 ; Cin = 1'b0 ; M = 1'b1 ;
#5; 
A = 4'b1100 ; B = 4'b1010 ; Cin = 1'b0 ; M = 1'b1 ;
#5; 
A = 4'b1100 ; B = 4'b1011 ; Cin = 1'b0 ; M = 1'b1 ;
#5; 
A = 4'b1100 ; B = 4'b1100 ; Cin = 1'b0 ; M = 1'b1 ;
#5; 
A = 4'b1100 ; B = 4'b1101 ; Cin = 1'b0 ; M = 1'b1 ;
#5; 
A = 4'b1100 ; B = 4'b1110 ; Cin = 1'b0 ; M = 1'b1 ;
#5; 
A = 4'b1100 ; B = 4'b1111 ; Cin = 1'b0 ; M = 1'b1 ;
#5; 
A = 4'b1101 ; B = 4'b0000 ; Cin = 1'b0 ; M = 1'b1 ;
#5; 
A = 4'b1101 ; B = 4'b0001 ; Cin = 1'b0 ; M = 1'b1 ;
#5; 
A = 4'b1101 ; B = 4'b0010 ; Cin = 1'b0 ; M = 1'b1 ;
#5; 
A = 4'b1101 ; B = 4'b0011 ; Cin = 1'b0 ; M = 1'b1 ;
#5; 
A = 4'b1101 ; B = 4'b0100 ; Cin = 1'b0 ; M = 1'b1 ;
#5; 
A = 4'b1101 ; B = 4'b0101 ; Cin = 1'b0 ; M = 1'b1 ;
#5; 
A = 4'b1101 ; B = 4'b0110 ; Cin = 1'b0 ; M = 1'b1 ;
#5; 
A = 4'b1101 ; B = 4'b0111 ; Cin = 1'b0 ; M = 1'b1 ;
#5; 
A = 4'b1101 ; B = 4'b1000 ; Cin = 1'b0 ; M = 1'b1 ;
#5; 
A = 4'b1101 ; B = 4'b1001 ; Cin = 1'b0 ; M = 1'b1 ;
#5; 
A = 4'b1101 ; B = 4'b1010 ; Cin = 1'b0 ; M = 1'b1 ;
#5; 
A = 4'b1101 ; B = 4'b1011 ; Cin = 1'b0 ; M = 1'b1 ;
#5; 
A = 4'b1101 ; B = 4'b1100 ; Cin = 1'b0 ; M = 1'b1 ;
#5; 
A = 4'b1101 ; B = 4'b1101 ; Cin = 1'b0 ; M = 1'b1 ;
#5; 
A = 4'b1101 ; B = 4'b1110 ; Cin = 1'b0 ; M = 1'b1 ;
#5; 
A = 4'b1101 ; B = 4'b1111 ; Cin = 1'b0 ; M = 1'b1 ;
#5; 
A = 4'b1110 ; B = 4'b0000 ; Cin = 1'b0 ; M = 1'b1 ;
#5; 
A = 4'b1110 ; B = 4'b0001 ; Cin = 1'b0 ; M = 1'b1 ;
#5; 
A = 4'b1110 ; B = 4'b0010 ; Cin = 1'b0 ; M = 1'b1 ;
#5; 
A = 4'b1110 ; B = 4'b0011 ; Cin = 1'b0 ; M = 1'b1 ;
#5; 
A = 4'b1110 ; B = 4'b0100 ; Cin = 1'b0 ; M = 1'b1 ;
#5; 
A = 4'b1110 ; B = 4'b0101 ; Cin = 1'b0 ; M = 1'b1 ;
#5; 
A = 4'b1110 ; B = 4'b0110 ; Cin = 1'b0 ; M = 1'b1 ;
#5; 
A = 4'b1110 ; B = 4'b0111 ; Cin = 1'b0 ; M = 1'b1 ;
#5; 
A = 4'b1110 ; B = 4'b1000 ; Cin = 1'b0 ; M = 1'b1 ;
#5; 
A = 4'b1110 ; B = 4'b1001 ; Cin = 1'b0 ; M = 1'b1 ;
#5; 
A = 4'b1110 ; B = 4'b1010 ; Cin = 1'b0 ; M = 1'b1 ;
#5; 
A = 4'b1110 ; B = 4'b1011 ; Cin = 1'b0 ; M = 1'b1 ;
#5; 
A = 4'b1110 ; B = 4'b1100 ; Cin = 1'b0 ; M = 1'b1 ;
#5; 
A = 4'b1110 ; B = 4'b1101 ; Cin = 1'b0 ; M = 1'b1 ;
#5; 
A = 4'b1110 ; B = 4'b1110 ; Cin = 1'b0 ; M = 1'b1 ;
#5; 
A = 4'b1110 ; B = 4'b1111 ; Cin = 1'b0 ; M = 1'b1 ;
#5; 
A = 4'b1111 ; B = 4'b0000 ; Cin = 1'b0 ; M = 1'b1 ;
#5; 
A = 4'b1111 ; B = 4'b0001 ; Cin = 1'b0 ; M = 1'b1 ;
#5; 
A = 4'b1111 ; B = 4'b0010 ; Cin = 1'b0 ; M = 1'b1 ;
#5; 
A = 4'b1111 ; B = 4'b0011 ; Cin = 1'b0 ; M = 1'b1 ;
#5; 
A = 4'b1111 ; B = 4'b0100 ; Cin = 1'b0 ; M = 1'b1 ;
#5; 
A = 4'b1111 ; B = 4'b0101 ; Cin = 1'b0 ; M = 1'b1 ;
#5; 
A = 4'b1111 ; B = 4'b0110 ; Cin = 1'b0 ; M = 1'b1 ;
#5; 
A = 4'b1111 ; B = 4'b0111 ; Cin = 1'b0 ; M = 1'b1 ;
#5; 
A = 4'b1111 ; B = 4'b1000 ; Cin = 1'b0 ; M = 1'b1 ;
#5; 
A = 4'b1111 ; B = 4'b1001 ; Cin = 1'b0 ; M = 1'b1 ;
#5; 
A = 4'b1111 ; B = 4'b1010 ; Cin = 1'b0 ; M = 1'b1 ;
#5; 
A = 4'b1111 ; B = 4'b1011 ; Cin = 1'b0 ; M = 1'b1 ;
#5; 
A = 4'b1111 ; B = 4'b1100 ; Cin = 1'b0 ; M = 1'b1 ;
#5; 
A = 4'b1111 ; B = 4'b1101 ; Cin = 1'b0 ; M = 1'b1 ;
#5; 
A = 4'b1111 ; B = 4'b1110 ; Cin = 1'b0 ; M = 1'b1 ;
#5; 
A = 4'b1111 ; B = 4'b1111 ; Cin = 1'b0 ; M = 1'b1 ;
#5; 
A = 4'b1111 ; B = 4'b1111 ; Cin = 1'b0 ; M = 1'b1 ;
end
endmodule



